module test_din#(
	parameter DWIDTH = 16
) (
	input clk,
	input rst_n,
	input din_valid,
	input [DWIDTH - 1 : 0] din_data
);

// work here

endmodule
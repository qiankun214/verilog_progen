module test_dout#(
	parameter DWIDTH = 16
) (
	input clk,
	input rst_n,
	output dout_valid,
	output [DWIDTH - 1 : 0] dout_data
);

// work here

endmodule
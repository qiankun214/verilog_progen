
// pro-gen:start here,coding before this line
module test_din #(
	parameter DWIDTH = 16
) (
	input rst_n,
	input din_valid,
	input clk,
	input [DWIDTH - 1 : 0] din_data
);

// link

// this on link:
	// 
// pro-gen:stop here,coding after this line
endmodule
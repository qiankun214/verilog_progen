// pro-gen:start here,coding before this line
module test_din#(
	parameter DWIDTH = 16
) (
	input rst_n,
	input din_valid,
	input [DWIDTH - 1 : 0] din_data,
	input clk
);


// pro-gen:stop here,coding after this line


endmodule
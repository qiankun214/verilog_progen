
// pro-gen:start here,coding before this line
module test_dout #(
	parameter DWIDTH = 16
) (
	input rst_n,
	output dout_valid,
	input clk,
	output [DWIDTH - 1 : 0] dout_data
);

// link

// this on link:
	// 
// pro-gen:stop here,coding after this line
endmodule
module test_dout#(
	parameter DWIDTH = 16
) (
	output [DWIDTH - 1 : 0] dout_data,
	output dout_valid,
	input rst_n,
	input clk
);

//progen-spilt:work after here


endmodule
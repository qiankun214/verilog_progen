module test_dout#(
	parameter DWIDTH = 16
) (
	input rst_n,
	output [DWIDTH - 1 : 0] dout_data,
	input clk,
	output dout_valid
);


//progen-spilt:work after here


endmodule
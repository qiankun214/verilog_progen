
// pro-gen:start here,coding before this line
module test_din #(
	parameter DWIDTH = 16
) (
	input clk,
	input rst_n,
	input din_valid,
	input [2 * DWIDTH + 3 - 1 : 0] din_data
);

// link

// this on link:
	// 
// pro-gen:stop here,coding after this line
endmodule
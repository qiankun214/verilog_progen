module test_din#(
	parameter DWIDTH = 16
) (
	input rst_n,
	input din_valid,
	input [DWIDTH - 1 : 0] din_data,
	input clk
);


//progen-spilt:work after here


endmodule
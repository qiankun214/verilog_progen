// pro-gen:start here,coding before this line
module test_dout#(
	parameter DWIDTH = 16
) (
	input rst_n,
	output [DWIDTH - 1 : 0] dout_data,
	input clk,
	output dout_valid
);


// pro-gen:stop here,coding after this line


endmodule
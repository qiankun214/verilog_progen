module test_din#(
	parameter DWIDTH = 16
) (
	input din_valid,
	input clk,
	input rst_n,
	input [DWIDTH - 1 : 0] din_data
);

None
// work here

endmodule